-------------------------------------------------------------------
--
--  Fichero:
--    rs232transmitter.vhd  15/7/2015
--
--    (c) J.M. Mendias
--    Dise�o Autom�tico de Sistemas
--    Facultad de Inform�tica. Universidad Complutense de Madrid
--
--  Prop�sito:
--    Conversor elemental de paralelo a una linea serie RS-232 con 
--    protocolo de strobe
--
--  Notas de dise�o:
--    - Parity: NONE
--    - Num data bits: 8
--    - Num stop bits: 1
--
-------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

entity rs232transmitter is
  generic (
    FREQ_KHZ : natural;  -- frecuencia de operacion en KHz
    BAUDRATE : natural   -- velocidad de comunicacion
  );
  port (
    -- host side
    clk     : in  std_logic;   -- reloj del sistema
    rst     : in  std_logic;   -- reset s�ncrono del sistema
    dataRdy : in  std_logic;   -- se activa durante 1 ciclo cada vez que hay un nuevo dato a transmitir
    data    : in  std_logic_vector (7 downto 0);   -- dato a transmitir
    busy    : out std_logic;   -- se activa mientras esta transmitiendo
    -- RS232 side
    TxD     : out std_logic    -- salida de datos serie del interfaz RS-232
  );
end rs232transmitter;

-------------------------------------------------------------------

use work.common.all;

architecture syn of rs232transmitter is

  signal baudCntCE, writeTxD : boolean;

begin

  baudCnt:
  process (clk)
    constant CYCLES : natural := (FREQ_KHZ*1000)/BAUDRATE;
    variable count  : natural range 0 to CYCLES-1 := 0;
  begin
    writeTxD <= (count = CYCLES-1);
    if rising_edge(clk) then
      if baudCntCE then
        count := (count + 1) mod CYCLES; 
      else
        count := 0;
      end if;
    end if;
  end process;
  
  fsmd:
  process (clk)
    variable bitPos : natural range 0 to 10 := 0;   
    variable TxDShf : std_logic_vector(9 downto 0) := (others =>'1');
  begin
    TxD <= TxDShf(0);
    --if baudCntCE then                         -- Esto esta mal ya que hace que busy dependa combinacionalmente de baudCntCE
    --  busy <= '1';                            -- Esto hace que se genere la señal con un ciclo de retraso, haciendo que
    --else                                      -- la fifo se desincronice
    --  busy <= '0';
    ---end if;
    if rising_edge(clk) then
      if rst='1' then
        TxDShf := (others =>'1'); 
        bitPos := 0;
      else
        case bitPos is
          when 0 =>                             -- Esperando solicitud de envio
            baudCntCE <= false;
            busy <= '0';                        -- Busy tiene que ser una señal moore 
            if dataRdy='1' then
              TxDShf := "1" & data & "0";
              bitPos := 1;
            end if;
          when others =>                        -- Desplaza
            baudCntCE <= true;
            busy <= '1';                        --Busy tiene que ser una señal moore 
            if writeTxD then
              TxDShf := "1" & TxDShf(9 downto 1);
              bitPos := (bitPos + 1) mod 11;
            end if;
        end case;
      end if;
    end if;
  end process;
  
end syn;

