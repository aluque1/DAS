LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY proyecto IS
  PORT (
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    ps2Clk : IN STD_LOGIC;
    ps2Data : IN STD_LOGIC;
    hSync : OUT STD_LOGIC;
    vSync : OUT STD_LOGIC;
    RGB : OUT STD_LOGIC_VECTOR(3 * 4 - 1 DOWNTO 0)
  );
END proyecto;

---------------------------------------------------------------------

LIBRARY ieee;
USE ieee.numeric_std.ALL;
USE work.common.ALL;

ARCHITECTURE syn OF proyecto IS

  CONSTANT FREQ_KHZ : NATURAL := 100_000; -- frecuencia de operacion en KHz
  CONSTANT VGA_KHZ : NATURAL := 25_000; -- frecuencia de envio de pixeles a la VGA en KHz
  CONSTANT FREQ_DIV : NATURAL := FREQ_KHZ/VGA_KHZ;
  constant negro : STD_LOGIC_VECTOR(11 DOWNTO 0) := "000000000000";
  constant grisOscuro : STD_LOGIC_VECTOR(11 DOWNTO 0) := "011101110111";
  constant grisClaro : STD_LOGIC_VECTOR(11 DOWNTO 0) := "100110011001";
  constant amarilloOscuro : STD_LOGIC_VECTOR(11 DOWNTO 0) := "110111010000";
  constant amarilloClaro : STD_LOGIC_VECTOR(11 DOWNTO 0) := "111111110000";
  constant azulOscuro : STD_LOGIC_VECTOR(11 DOWNTO 0) := "";
  constant azulClaro : STD_LOGIC_VECTOR(11 DOWNTO 0) := "";
  
  signal xPiezaAct : unsigned(7 downto 0) := to_unsigned(5, 8);
  signal yPiezaAct : unsigned(7 downto 0) := to_unsigned(0, 8);
  
  signal addrTabRd : unsigned(7 downto 0) := (others => '0');
  signal addrTabWr : unsigned(7 downto 0) := (others => '0');
  
  signal distASuelo : natural := 2; -- variable que se modifica
  
  SIGNAL aP, sP, dP, rP, spcP, actCuadrado, actLinea, lineaPos1, lineaPos2 : BOOLEAN := false;

  SIGNAL rstSync : STD_LOGIC;
  SIGNAL data : STD_LOGIC_VECTOR(7 DOWNTO 0);
  SIGNAL dataRdy : STD_LOGIC;

  SIGNAL color : STD_LOGIC_VECTOR(11 DOWNTO 0);
  signal colorPiezaActB : std_logic_vector (11 downto 0) := amarilloClaro;
  signal colorPiezaActI : std_logic_vector (11 downto 0) := amarilloOscuro;
  
  signal visual: std_logic_vector(3 downto 0) := (others => '0');--Muy seguramente aumenten los bits
  --visual(0) bordes claritos de los bordes del campo
  --visual(1) interior oscuro
  --visual(2) lineas de las piezas
  --visual(3) relleno de las piezas
  --A IMPLEMENTAR
  --visual(4) lineas piezas en el campo
  --visual(5) relleno piezas en el campo
  SIGNAL cuadradoB, cuadradoI, piezaActualB, piezaActualI: STD_LOGIC;
  SIGNAL mover, finPartida, reiniciar : BOOLEAN;

  type tablero_t is array (0 to 230) of unsigned(2 downto 0); 
  signal tablero : tablero_t := (others => (others => '0'));

  SIGNAL lineAux, pixelAux : STD_LOGIC_VECTOR(9 DOWNTO 0);
  SIGNAL line, pixel : unsigned(7 DOWNTO 0);
  
  signal x : natural := 14;
  signal y : natural := 54;
  
BEGIN

  rstSynchronizer : synchronizer
  GENERIC MAP(STAGES => 2, XPOL => '0')
  PORT MAP(clk => clk, x => rst, xSync => rstSync);

  ------------------  

  ps2KeyboardInterface : ps2receiver
  PORT MAP(clk => clk, rst => rstSync, dataRdy => dataRdy, data => data, ps2Clk => ps2Clk, ps2Data => ps2Data);

  keyboardScanner :
  PROCESS (clk)
    TYPE states IS (keyON, keyOFF);
    VARIABLE state : states := keyON; --Puede estar mal no se
  BEGIN
    IF rising_edge(clk) THEN
      IF rstSync = '1' THEN
        state := keyOFF; --Revisar lo de el estado inicial
      ELSIF dataRdy = '1' THEN
        CASE state IS
          WHEN keyON =>
            CASE data IS
              WHEN X"F0" => state := keyOFF;
              WHEN X"1C" => aP <= true;
              WHEN X"1B" => sP <= true;
              WHEN X"23" => dP <= true;
              WHEN X"2D" => rP <= true;
              WHEN X"29" => spcP <= true;
              WHEN OTHERS => state := keyON;
            END CASE;
          WHEN keyOFF =>
            state := keyON;
            CASE data IS
              WHEN X"1C" => aP <= false;
              WHEN X"1B" => sP <= false;
              WHEN X"23" => dP <= false;
              WHEN X"2D" => rP <= false;
              WHEN X"29" => spcP <= false;
              WHEN OTHERS => state := keyOFF;
            END CASE;
        END CASE;
      END IF;
    END IF;
  END PROCESS;

  ------------------  

  screenInteface : vgaRefresher
  GENERIC MAP(FREQ_DIV => FREQ_DIV)
  PORT MAP(clk => clk, line => lineAux, pixel => pixelAux, R => color(11 downto 8), G => color(7 downto 4), B => color(3 downto 0), hSync => hSync, vSync => vSync, RGB => RGB);

  pixel <= unsigned(pixelAux(9 DOWNTO 2));
  line <= unsigned(lineAux(9 DOWNTO 2));

  with visual select
    color <= 
    grisClaro when "0001",
    grisOscuro when "0010",
    grisClaro when "0011",
    colorPiezaActB when "0100",
    colorPiezaActB when "1100",
    colorPiezaActI when "1000",
    negro when others;
    
  ------------------

  
  visual(0) <= '1' when (pixel = y and ((line > 9 and line < 14) or (line > 114 and line < 119))) or
                        (line = x and ((pixel > 49 and pixel < 54) or (pixel > 104 and pixel < 109))) or
                        (line = 9 and (pixel >= 49 and pixel <= 109)) or
                        (line = 14 and (pixel >= 54 and pixel <= 104)) or
                        (line = 114 and (pixel >= 54 and pixel <= 104)) or
                        (line = 119 and (pixel >= 49 and pixel <= 109)) or
                        (pixel = 49 and (line >= 9 and line <= 119)) or
                        (pixel = 54 and (line >= 14 and line <= 114)) or
                        (pixel = 104 and (line >= 14 and line <= 114)) or
                        (pixel = 109 and (line >= 9 and line <= 119)) else '0';
                        
  visual(1) <= '1' when ((pixel > 49 and pixel < 109) and ((line > 9 and line < 14) or (line > 114 and line < 119))) or
                        ((line > 9 and line < 119) and ((pixel > 49 and pixel < 54) or (pixel > 104 and pixel < 109))) else '0';
  
  visual(2) <= '1' when piezaActualB = '1' else '0';
  
  visual(3) <= '1' when piezaActualI = '1' else '0';
  
  piezaActualB <= '1' when cuadradoB = '1' else '0'; --piezaActualB <= '1' when cuadradoB = '1' or .... else '0';
  piezaActualI <= '1' when cuadradoI = '1' else '0'; --piezaActualI <= '1' when cuadradoI = '1' or .... else '0';
  
  cuadradoB <= '1' when ((pixel = xPiezaAct or pixel = (xPiezaAct + 10) or pixel = (xPiezaAct + 5)) and (line >= yPiezaAct and line <= (yPiezaAct + 10))) or
                         ((line = yPiezaAct or line = (yPiezaAct + 10) or line = (yPiezaAct + 5)) and (pixel >= xPiezaAct and pixel <= (xPiezaAct + 10))) else '0';
                         --Aqui poner variable que le indique cuando pintarse
  cuadradoI <= '1' when (pixel > xPiezaAct and pixel < (xPiezaAct + 10)) and (line > yPiezaAct and line < (yPiezaAct + 10)) else '0';
  
  pulseGen :
  PROCESS (clk)
    CONSTANT CYCLES : NATURAL := hz2cycles(FREQ_KHZ, 50);
    VARIABLE count : NATURAL RANGE 0 TO CYCLES - 1 := 0;
  BEGIN
    IF rising_edge(clk) THEN
      IF rstSync = '1' THEN
        count := 0;
      ELSIF finPartida = false THEN
        count := (count + 1) MOD CYCLES;
        mover <= false;
        IF count = (CYCLES - 1) THEN
          mover <= true;
        END IF;
      END IF;
    END IF;
  END PROCESS;

  ------------------
  --Replantear el movimiento entero de la pieza
  movPiezaTab:
  process(clk)
  begin
    if rising_edge(clk) then
        if mover then
            if yPiezaAct + distASuelo < 220 and ... and (xPiezaAct > 0 and xPiezaAct < 11) then --falta la se�al colision
                --Aqui se manda la se�al para borrar la pieza
                if sP then
                    yPiezaAct <= yPiezaAct + 2;
                else
                    yPiezaAct <= yPiezaAct + 1;
                end if;
                if aP then
                    xPiezaAct <= xPiezaAct - 1;
                end if;
                if dP then
                    xPiezaAct <= xPiezaAct + 1;
                end if;
            end if;
        end if;
    end if;
  end process;


  ------------------

 
  regSumX:
  process(clk)
  begin
    if rising_edge(clk) then
        if (line = x+1 and ((pixel > 49 and pixel < 54) or (pixel > 104 and pixel < 109))) then
            x <= x + 5;
            if x = 114 then
                x <= 14;
            end if;
        end if;
    end if;
  end process;
  
  regSumY:
  process(clk)
  begin
  if rising_edge(clk) then
        if (pixel = y+1 and ((line > 9 and line < 14) or (line > 114 and line < 119))) then
            y <= y + 5;
            if y = 104 then
                y <= 54;
            end if;
        end if;
    end if;
  end process;

-------------------------------------------
--Limpiado, dibujado de piezas y colision--
-------------------------------------------
--Falta implementar lo de colision
--A lo mejor hay que meter una se�al para mandar el limpiado a la hora de darle a la r
---------------------------------
  limpiaCuadrado:
  tablero(to_integer(11*yPiezaAct + xPiezaAct)) <= (others => '0') when actCuadrado else tablero(to_integer(11*yPiezaAct + xPiezaAct));
  tablero(to_integer(11*yPiezaAct + (xPiezaAct+1))) <= (others => '0') when actCuadrado else tablero(to_integer(11*yPiezaAct + (xPiezaAct+1)));
  tablero(to_integer(11*(yPiezaAct+1) + xPiezaAct)) <= (others => '0') when actCuadrado else tablero(to_integer(11*(yPiezaAct+1) + xPiezaAct));
  tablero(to_integer(11*(yPiezaAct+1) + (xPiezaAct+1))) <= (others => '0') when actCuadrado else tablero(to_integer(11*(yPiezaAct+1) + (xPiezaAct+1)));
  
  pintaCuadrado:
  tablero(to_integer(11*yPiezaAct + xPiezaAct)) <= to_unsigned(1,3) when actCuadrado else tablero(to_integer(11*yPiezaAct + xPiezaAct));
  tablero(to_integer(11*yPiezaAct + (xPiezaAct+1))) <= to_unsigned(1,3) when actCuadrado else tablero(to_integer(11*yPiezaAct + (xPiezaAct+1)));
  tablero(to_integer(11*(yPiezaAct+1) + xPiezaAct)) <= to_unsigned(1,3) when actCuadrado else tablero(to_integer(11*(yPiezaAct+1) + xPiezaAct));
  tablero(to_integer(11*(yPiezaAct+1) + (xPiezaAct+1))) <= to_unsigned(1,3) when actCuadrado else tablero(to_integer(11*(yPiezaAct+1) + (xPiezaAct+1)));
  
---------------------------------
   
  limpiaLineaPos1:
  tablero(to_integer(11*yPiezaAct + xPiezaAct)) <= (others => '0') when actLinea and lineaPos1 else tablero(to_integer(11*yPiezaAct + xPiezaAct));
  tablero(to_integer(11*yPiezaAct + (xPiezaAct+1))) <= (others => '0') when actLinea and lineaPos1 else tablero(to_integer(11*yPiezaAct + (xPiezaAct+1)));
  tablero(to_integer(11*yPiezaAct + (xPiezaAct+2))) <= (others => '0') when actLinea and lineaPos1 else tablero(to_integer(11*yPiezaAct + (xPiezaAct+2)));
  tablero(to_integer(11*yPiezaAct + (xPiezaAct+3))) <= (others => '0') when actLinea and lineaPos1 else tablero(to_integer(11*yPiezaAct + (xPiezaAct+3)));
  
  pintaLineaPos1:
  tablero(to_integer(11*yPiezaAct + xPiezaAct)) <= to_unsigned(2,3) when actLinea and lineaPos1 else tablero(to_integer(11*yPiezaAct + xPiezaAct));
  tablero(to_integer(11*yPiezaAct + (xPiezaAct+1))) <= to_unsigned(2,3) when actLinea and lineaPos1 else tablero(to_integer(11*yPiezaAct + (xPiezaAct+1)));
  tablero(to_integer(11*yPiezaAct + (xPiezaAct+2))) <= to_unsigned(2,3) when actLinea and lineaPos1 else tablero(to_integer(11*yPiezaAct + (xPiezaAct+2)));
  tablero(to_integer(11*yPiezaAct + (xPiezaAct+3))) <= to_unsigned(2,3) when actLinea and lineaPos1 else tablero(to_integer(11*yPiezaAct + (xPiezaAct+3)));
  
  limpiaLineaPos2:
  tablero(to_integer(11*yPiezaAct + xPiezaAct)) <= (others => '0') when actLinea and lineaPos2 else tablero(to_integer(11*yPiezaAct + xPiezaAct));
  tablero(to_integer(11*(yPiezaAct+1) + xPiezaAct)) <= (others => '0') when actLinea and lineaPos2 else tablero(to_integer(11*(yPiezaAct+1) + xPiezaAct));
  tablero(to_integer(11*(yPiezaAct+2) + xPiezaAct)) <= (others => '0') when actLinea and lineaPos2 else tablero(to_integer(11*(yPiezaAct+2) + xPiezaAct));
  tablero(to_integer(11*(yPiezaAct+3) + xPiezaAct)) <= (others => '0') when actLinea and lineaPos2 else tablero(to_integer(11*(yPiezaAct+3) + xPiezaAct));
  
  pintaLineaPos2:
  tablero(to_integer(11*yPiezaAct + xPiezaAct)) <= to_unsigned(2,3) when actLinea and lineaPos2 else tablero(to_integer(11*yPiezaAct + xPiezaAct));
  tablero(to_integer(11*(yPiezaAct+1) + xPiezaAct)) <= to_unsigned(2,3) when actLinea and lineaPos2 else tablero(to_integer(11*(yPiezaAct+1) + xPiezaAct));
  tablero(to_integer(11*(yPiezaAct+2) + xPiezaAct)) <= to_unsigned(2,3) when actLinea and lineaPos2 else tablero(to_integer(11*(yPiezaAct+2) + xPiezaAct));
  tablero(to_integer(11*(yPiezaAct+3) + xPiezaAct)) <= to_unsigned(2,3) when actLinea and lineaPos2 else tablero(to_integer(11*(yPiezaAct+3) + xPiezaAct));

---------------------------------

  limpiaZetaPos1:
  tablero(to_integer(11*yPiezaAct + xPiezaAct)) <= (others => '0') when ... else tablero(to_integer(11*yPiezaAct + xPiezaAct));
  tablero(to_integer(11*yPiezaAct + (xPiezaAct+1))) <= (others => '0') when ... else tablero(to_integer(11*yPiezaAct + (xPiezaAct+1)));
  tablero(to_integer(11*(yPiezaAct+1) + (xPiezaAct+1))) <= (others => '0') when ... else tablero(to_integer(11*(yPiezaAct+1) + (xPiezaAct+1)));
  tablero(to_integer(11*(yPiezaAct+2) + (xPiezaAct+1))) <= (others => '0') when ... else tablero(to_integer(11*(yPiezaAct+2) + (xPiezaAct+1)));
  tablero(to_integer(11*(yPiezaAct+2) + (xPiezaAct+2))) <= (others => '0') when ... else tablero(to_integer(11*(yPiezaAct+2) + (xPiezaAct+2)));
  
  pintaZetaPos1:
  tablero(to_integer(11*yPiezaAct + xPiezaAct)) <= to_unsigned(3,3) when ... else tablero(to_integer(11*yPiezaAct + xPiezaAct));
  tablero(to_integer(11*yPiezaAct + (xPiezaAct+1))) <= to_unsigned(3,3) when ... else tablero(to_integer(11*yPiezaAct + (xPiezaAct+1)));
  tablero(to_integer(11*(yPiezaAct+1) + (xPiezaAct+1))) <= to_unsigned(3,3) when ... else tablero(to_integer(11*(yPiezaAct+1) + (xPiezaAct+1)));
  tablero(to_integer(11*(yPiezaAct+2) + (xPiezaAct+1))) <= to_unsigned(3,3) when ... else tablero(to_integer(11*(yPiezaAct+2) + (xPiezaAct+1)));
  tablero(to_integer(11*(yPiezaAct+2) + (xPiezaAct+2))) <= to_unsigned(3,3) when ... else tablero(to_integer(11*(yPiezaAct+2) + (xPiezaAct+2)));
  
  limpiaZetaPos2:
  tablero(to_integer(11*yPiezaAct + xPiezaAct)) <= (others => '0') when ... else tablero(to_integer(11*yPiezaAct + xPiezaAct));
  tablero(to_integer(11*(yPiezaAct+1) + xPiezaAct)) <= (others => '0') when ... else tablero(to_integer(11*(yPiezaAct+1) + xPiezaAct));
  tablero(to_integer(11*yPiezaAct + (xPiezaAct+1))) <= (others => '0') when ... else tablero(to_integer(11*yPiezaAct + (xPiezaAct+1)));
  tablero(to_integer(11*yPiezaAct + (xPiezaAct+2))) <= (others => '0') when ... else tablero(to_integer(11*yPiezaAct + (xPiezaAct+2)));
  tablero(to_integer(11*(yPiezaAct-1) + (xPiezaAct+2))) <= (others => '0') when ... else tablero(to_integer(11*(yPiezaAct-1) + (xPiezaAct+2)));
  
  pintaZetaPos2:
  tablero(to_integer(11*yPiezaAct + xPiezaAct)) <= to_unsigned(3,3) when ... else tablero(to_integer(11*yPiezaAct + xPiezaAct));
  tablero(to_integer(11*(yPiezaAct+1) + xPiezaAct)) <= to_unsigned(3,3) when ... else tablero(to_integer(11*(yPiezaAct+1) + xPiezaAct));
  tablero(to_integer(11*yPiezaAct + (xPiezaAct+1))) <= to_unsigned(3,3) when ... else tablero(to_integer(11*yPiezaAct + (xPiezaAct+1)));
  tablero(to_integer(11*yPiezaAct + (xPiezaAct+2))) <= to_unsigned(3,3) when ... else tablero(to_integer(11*yPiezaAct + (xPiezaAct+2)));
  tablero(to_integer(11*(yPiezaAct-1) + (xPiezaAct+2))) <= to_unsigned(3,3) when ... else tablero(to_integer(11*(yPiezaAct-1) + (xPiezaAct+2)));
  
---------------------------------
  
  limpiaZetaInvPos1:
  tablero(to_integer(11*yPiezaAct + xPiezaAct)) <= (others => '0') when ... else tablero(to_integer(11*yPiezaAct + xPiezaAct));
  tablero(to_integer(11*yPiezaAct + (xPiezaAct+1))) <= (others => '0') when ... else tablero(to_integer(11*yPiezaAct + (xPiezaAct+1)));
  tablero(to_integer(11*(yPiezaAct+1) + xPiezaAct)) <= (others => '0') when ... else tablero(to_integer(11*(yPiezaAct+1) + xPiezaAct));
  tablero(to_integer(11*(yPiezaAct+2) + xPiezaAct)) <= (others => '0') when ... else tablero(to_integer(11*(yPiezaAct+2) + xPiezaAct));
  tablero(to_integer(11*(yPiezaAct+2) + (xPiezaAct-1))) <= (others => '0') when ... else tablero(to_integer(11*(yPiezaAct+2) + (xPiezaAct-1)));
  
  pintaZetaInvPos1:
  tablero(to_integer(11*yPiezaAct + xPiezaAct)) <= to_unsigned(4,3) when ... else tablero(to_integer(11*yPiezaAct + xPiezaAct));
  tablero(to_integer(11*yPiezaAct + (xPiezaAct+1))) <= to_unsigned(4,3) when ... else tablero(to_integer(11*yPiezaAct + (xPiezaAct+1)));
  tablero(to_integer(11*(yPiezaAct+1) + xPiezaAct)) <= to_unsigned(4,3) when ... else tablero(to_integer(11*(yPiezaAct+1) + xPiezaAct));
  tablero(to_integer(11*(yPiezaAct+2) + xPiezaAct)) <= to_unsigned(4,3) when ... else tablero(to_integer(11*(yPiezaAct+2) + xPiezaAct));
  tablero(to_integer(11*(yPiezaAct+2) + (xPiezaAct-1))) <= to_unsigned(4,3) when ... else tablero(to_integer(11*(yPiezaAct+2) + (xPiezaAct-1)));
  
  limpiaZetaInvPos2:
  tablero(to_integer(11*yPiezaAct + xPiezaAct)) <= (others => '0') when ... else tablero(to_integer(11*yPiezaAct + xPiezaAct));
  tablero(to_integer(11*(yPiezaAct+1) + xPiezaAct)) <= (others => '0') when ... else tablero(to_integer(11*(yPiezaAct+1) + xPiezaAct));
  tablero(to_integer(11*(yPiezaAct+1) + (xPiezaAct+1))) <= (others => '0') when ... else tablero(to_integer(11*(yPiezaAct+1) + (xPiezaAct+1)));
  tablero(to_integer(11*(yPiezaAct+1) + (xPiezaAct+2))) <= (others => '0') when ... else tablero(to_integer(11*(yPiezaAct+1) + (xPiezaAct+2)));
  tablero(to_integer(11*(yPiezaAct+2) + (xPiezaAct+2))) <= (others => '0') when ... else tablero(to_integer(11*(yPiezaAct+2) + (xPiezaAct+2)));
  
  pintaZetaInvPos2:
  tablero(to_integer(11*yPiezaAct + xPiezaAct)) <= to_unsigned(4,3) when ... else tablero(to_integer(11*yPiezaAct + xPiezaAct));
  tablero(to_integer(11*(yPiezaAct+1) + xPiezaAct)) <= to_unsigned(4,3) when ... else tablero(to_integer(11*(yPiezaAct+1) + xPiezaAct));
  tablero(to_integer(11*(yPiezaAct+1) + (xPiezaAct+1))) <= to_unsigned(4,3) when ... else tablero(to_integer(11*(yPiezaAct+1) + (xPiezaAct+1)));
  tablero(to_integer(11*(yPiezaAct+1) + (xPiezaAct+2))) <= to_unsigned(4,3) when ... else tablero(to_integer(11*(yPiezaAct+1) + (xPiezaAct+2)));
  tablero(to_integer(11*(yPiezaAct+2) + (xPiezaAct+2))) <= to_unsigned(4,3) when ... else tablero(to_integer(11*(yPiezaAct+2) + (xPiezaAct+2)));
  
---------------------------------
  
  limpiaElePos1:
  tablero(to_integer(11*yPiezaAct + xPiezaAct)) <= (others => '0') when ... else tablero(to_integer(11*yPiezaAct + xPiezaAct));
  tablero(to_integer(11*(yPiezaAct+1) + xPiezaAct)) <= (others => '0') when ... else tablero(to_integer(11*(yPiezaAct+1) + xPiezaAct));
  tablero(to_integer(11*(yPiezaAct+2) + xPiezaAct)) <= (others => '0') when ... else tablero(to_integer(11*(yPiezaAct+2) + xPiezaAct));
  tablero(to_integer(11*(yPiezaAct+2) + (xPiezaAct+1))) <= (others => '0') when ... else tablero(to_integer(11*(yPiezaAct+2) + (xPiezaAct+1)));
  
  pintaElePos1:
  tablero(to_integer(11*yPiezaAct + xPiezaAct)) <= to_unsigned(5,3) when ... else tablero(to_integer(11*yPiezaAct + xPiezaAct));
  tablero(to_integer(11*(yPiezaAct+1) + xPiezaAct)) <= to_unsigned(5,3) when ... else tablero(to_integer(11*(yPiezaAct+1) + xPiezaAct));
  tablero(to_integer(11*(yPiezaAct+2) + xPiezaAct)) <= to_unsigned(5,3) when ... else tablero(to_integer(11*(yPiezaAct+2) + xPiezaAct));
  tablero(to_integer(11*(yPiezaAct+2) + (xPiezaAct+1))) <= to_unsigned(5,3) when ... else tablero(to_integer(11*(yPiezaAct+2) + (xPiezaAct+1)));
  
  limpiaElePos2:
  tablero(to_integer(11*yPiezaAct + xPiezaAct)) <= (others => '0') when ... else tablero(to_integer(11*yPiezaAct + xPiezaAct));
  tablero(to_integer(11*(yPiezaAct+1) + xPiezaAct)) <= (others => '0') when ... else tablero(to_integer(11*(yPiezaAct+1) + xPiezaAct));
  tablero(to_integer(11*yPiezaAct + (xPiezaAct+1))) <= (others => '0') when ... else tablero(to_integer(11*yPiezaAct + (xPiezaAct+1)));
  tablero(to_integer(11*yPiezaAct + (xPiezaAct+2))) <= (others => '0') when ... else tablero(to_integer(11*yPiezaAct + (xPiezaAct+2)));
  
  pintaElePos2:
  tablero(to_integer(11*yPiezaAct + xPiezaAct)) <= to_unsigned(5,3) when ... else tablero(to_integer(11*yPiezaAct + xPiezaAct));
  tablero(to_integer(11*(yPiezaAct+1) + xPiezaAct)) <= to_unsigned(5,3) when ... else tablero(to_integer(11*(yPiezaAct+1) + xPiezaAct));
  tablero(to_integer(11*yPiezaAct + (xPiezaAct+1))) <= to_unsigned(5,3) when ... else tablero(to_integer(11*yPiezaAct + (xPiezaAct+1)));
  tablero(to_integer(11*yPiezaAct + (xPiezaAct+2))) <= to_unsigned(5,3) when ... else tablero(to_integer(11*yPiezaAct + (xPiezaAct+2)));
  
  limpiaElePos3:
  tablero(to_integer(11*yPiezaAct + xPiezaAct)) <= (others => '0') when ... else tablero(to_integer(11*yPiezaAct + xPiezaAct));
  tablero(to_integer(11*yPiezaAct + (xPiezaAct+1))) <= (others => '0') when ... else tablero(to_integer(11*yPiezaAct + (xPiezaAct+1)));
  tablero(to_integer(11*(yPiezaAct+2) + (xPiezaAct+1))) <= (others => '0') when ... else tablero(to_integer(11*(yPiezaAct+2) + (xPiezaAct+1)));
  tablero(to_integer(11*(yPiezaAct+3) + (xPiezaAct+1))) <= (others => '0') when ... else tablero(to_integer(11*(yPiezaAct+3) + (xPiezaAct+1)));
   
  pintaElePos3:
  tablero(to_integer(11*yPiezaAct + xPiezaAct)) <= to_unsigned(5,3) when ... else tablero(to_integer(11*yPiezaAct + xPiezaAct));
  tablero(to_integer(11*yPiezaAct + (xPiezaAct+1))) <= to_unsigned(5,3) when ... else tablero(to_integer(11*yPiezaAct + (xPiezaAct+1)));
  tablero(to_integer(11*(yPiezaAct+2) + (xPiezaAct+1))) <= to_unsigned(5,3) when ... else tablero(to_integer(11*(yPiezaAct+2) + (xPiezaAct+1)));
  tablero(to_integer(11*(yPiezaAct+3) + (xPiezaAct+1))) <= to_unsigned(5,3) when ... else tablero(to_integer(11*(yPiezaAct+3) + (xPiezaAct+1)));
  
  limpiaElePos4:
  tablero(to_integer(11*yPiezaAct + xPiezaAct)) <= (others => '0') when ... else tablero(to_integer(11*yPiezaAct + xPiezaAct));
  tablero(to_integer(11*yPiezaAct + (xPiezaAct+1))) <= (others => '0') when ... else tablero(to_integer(11*yPiezaAct + (xPiezaAct+1)));
  tablero(to_integer(11*yPiezaAct + (xPiezaAct+2))) <= (others => '0') when ... else tablero(to_integer(11*yPiezaAct + (xPiezaAct+2)));
  tablero(to_integer(11*(yPiezaAct-1) + (xPiezaAct+2))) <= (others => '0') when ... else tablero(to_integer(11*(yPiezaAct-1) + (xPiezaAct+2)));
  
  pintaElePos4:
  tablero(to_integer(11*yPiezaAct + xPiezaAct)) <= to_unsigned(5,3) when ... else tablero(to_integer(11*yPiezaAct + xPiezaAct));
  tablero(to_integer(11*yPiezaAct + (xPiezaAct+1))) <= to_unsigned(5,3) when ... else tablero(to_integer(11*yPiezaAct + (xPiezaAct+1)));
  tablero(to_integer(11*yPiezaAct + (xPiezaAct+2))) <= to_unsigned(5,3) when ... else tablero(to_integer(11*yPiezaAct + (xPiezaAct+2)));
  tablero(to_integer(11*(yPiezaAct-1) + (xPiezaAct+2))) <= to_unsigned(5,3) when ... else tablero(to_integer(11*(yPiezaAct-1) + (xPiezaAct+2)));
  
---------------------------------
  
  limpiaEleInvPos1:
  tablero(to_integer(11*yPiezaAct + xPiezaAct)) <= (others => '0') when ... else tablero(to_integer(11*yPiezaAct + xPiezaAct));
  tablero(to_integer(11*(yPiezaAct+1) + xPiezaAct)) <= (others => '0') when ... else tablero(to_integer(11*(yPiezaAct+1) + xPiezaAct));
  tablero(to_integer(11*(yPiezaAct+2) + xPiezaAct)) <= (others => '0') when ... else tablero(to_integer(11*(yPiezaAct+2) + xPiezaAct));
  tablero(to_integer(11*(yPiezaAct+2) + (xPiezaAct-1))) <= (others => '0') when ... else tablero(to_integer(11*(yPiezaAct+2) + (xPiezaAct-1)));
  
  pintaEleInvPos1:
  tablero(to_integer(11*yPiezaAct + xPiezaAct)) <= to_unsigned(6,3) when ... else tablero(to_integer(11*yPiezaAct + xPiezaAct));
  tablero(to_integer(11*(yPiezaAct+1) + xPiezaAct)) <= to_unsigned(6,3) when ... else tablero(to_integer(11*(yPiezaAct+1) + xPiezaAct));
  tablero(to_integer(11*(yPiezaAct+2) + xPiezaAct)) <= to_unsigned(6,3) when ... else tablero(to_integer(11*(yPiezaAct+2) + xPiezaAct));
  tablero(to_integer(11*(yPiezaAct+2) + (xPiezaAct-1))) <= to_unsigned(6,3) when ... else tablero(to_integer(11*(yPiezaAct+2) + (xPiezaAct-1)));
  
  limpiaEleInvPos2:
  tablero(to_integer(11*yPiezaAct + xPiezaAct)) <= (others => '0') when ... else tablero(to_integer(11*yPiezaAct + xPiezaAct));
  tablero(to_integer(11*(yPiezaAct+1) + xPiezaAct)) <= (others => '0') when ... else tablero(to_integer(11*(yPiezaAct+1) + xPiezaAct));
  tablero(to_integer(11*(yPiezaAct+1) + (xPiezaAct+1))) <= (others => '0') when ... else tablero(to_integer(11*(yPiezaAct+1) + (xPiezaAct+1)));
  tablero(to_integer(11*(yPiezaAct+1) + (xPiezaAct+2))) <= (others => '0') when ... else tablero(to_integer(11*(yPiezaAct+1) + (xPiezaAct+2)));
  
  pintaEleInvPos2:
  tablero(to_integer(11*yPiezaAct + xPiezaAct)) <= to_unsigned(6,3) when ... else tablero(to_integer(11*yPiezaAct + xPiezaAct));
  tablero(to_integer(11*(yPiezaAct+1) + xPiezaAct)) <= to_unsigned(6,3) when ... else tablero(to_integer(11*(yPiezaAct+1) + xPiezaAct));
  tablero(to_integer(11*(yPiezaAct+1) + (xPiezaAct+1))) <= to_unsigned(6,3) when ... else tablero(to_integer(11*(yPiezaAct+1) + (xPiezaAct+1)));
  tablero(to_integer(11*(yPiezaAct+1) + (xPiezaAct+2))) <= to_unsigned(6,3) when ... else tablero(to_integer(11*(yPiezaAct+1) + (xPiezaAct+2)));
  
  limpiaEleInvPos3:
  tablero(to_integer(11*yPiezaAct + xPiezaAct)) <= (others => '0') when ... else tablero(to_integer(11*yPiezaAct + xPiezaAct));
  tablero(to_integer(11*yPiezaAct + (xPiezaAct+1))) <= (others => '0') when ... else tablero(to_integer(11*yPiezaAct + (xPiezaAct+1)));
  tablero(to_integer(11*(yPiezaAct+2) + xPiezaAct)) <= (others => '0') when ... else tablero(to_integer(11*(yPiezaAct+2) + xPiezaAct));
  tablero(to_integer(11*(yPiezaAct+3) + xPiezaAct)) <= (others => '0') when ... else tablero(to_integer(11*(yPiezaAct+3) + xPiezaAct));
  
  pintaEleInvPos3:
  tablero(to_integer(11*yPiezaAct + xPiezaAct)) <= to_unsigned(6,3) when ... else tablero(to_integer(11*yPiezaAct + xPiezaAct));
  tablero(to_integer(11*yPiezaAct + (xPiezaAct+1))) <= to_unsigned(6,3) when ... else tablero(to_integer(11*yPiezaAct + (xPiezaAct+1)));
  tablero(to_integer(11*(yPiezaAct+2) + xPiezaAct)) <= to_unsigned(6,3) when ... else tablero(to_integer(11*(yPiezaAct+2) + xPiezaAct));
  tablero(to_integer(11*(yPiezaAct+3) + xPiezaAct)) <= to_unsigned(6,3) when ... else tablero(to_integer(11*(yPiezaAct+3) + xPiezaAct));
  
  limpiaEleInvPos4:
  tablero(to_integer(11*yPiezaAct + xPiezaAct)) <= (others => '0') when ... else tablero(to_integer(11*yPiezaAct + xPiezaAct));
  tablero(to_integer(11*yPiezaAct + (xPiezaAct+1))) <= (others => '0') when ... else tablero(to_integer(11*yPiezaAct + (xPiezaAct+1)));
  tablero(to_integer(11*yPiezaAct + (xPiezaAct+2))) <= (others => '0') when ... else tablero(to_integer(11*yPiezaAct + (xPiezaAct+2)));
  tablero(to_integer(11*(yPiezaAct+1) + (xPiezaAct+2))) <= (others => '0') when ... else tablero(to_integer(11*(yPiezaAct+1) + (xPiezaAct+2)));
  
  limpiaEleInvPos4:
  tablero(to_integer(11*yPiezaAct + xPiezaAct)) <= to_unsigned(6,3) when ... else tablero(to_integer(11*yPiezaAct + xPiezaAct));
  tablero(to_integer(11*yPiezaAct + (xPiezaAct+1))) <= to_unsigned(6,3) when ... else tablero(to_integer(11*yPiezaAct + (xPiezaAct+1)));
  tablero(to_integer(11*yPiezaAct + (xPiezaAct+2))) <= to_unsigned(6,3) when ... else tablero(to_integer(11*yPiezaAct + (xPiezaAct+2)));
  tablero(to_integer(11*(yPiezaAct+1) + (xPiezaAct+2))) <= to_unsigned(6,3) when ... else tablero(to_integer(11*(yPiezaAct+1) + (xPiezaAct+2)));
  
---------------------------------
  
  limpiaTePos1:
  tablero(to_integer(11*yPiezaAct + xPiezaAct)) <= (others => '0') when ... else tablero(to_integer(11*yPiezaAct + xPiezaAct));
  tablero(to_integer(11*(yPiezaAct+1) + xPiezaAct)) <= (others => '0') when ... else tablero(to_integer(11*(yPiezaAct+1) + xPiezaAct));
  tablero(to_integer(11*(yPiezaAct+2) + xPiezaAct)) <= (others => '0') when ... else tablero(to_integer(11*(yPiezaAct+2) + xPiezaAct));
  tablero(to_integer(11*(yPiezaAct+1) + (xPiezaAct-1))) <= (others => '0') when ... else tablero(to_integer(11*(yPiezaAct+1) + (xPiezaAct-1)));
   
  pintaTePos1:
  tablero(to_integer(11*yPiezaAct + xPiezaAct)) <= to_unsigned(7,3) when ... else tablero(to_integer(11*yPiezaAct + xPiezaAct));
  tablero(to_integer(11*(yPiezaAct+1) + xPiezaAct)) <= to_unsigned(7,3) when ... else tablero(to_integer(11*(yPiezaAct+1) + xPiezaAct));
  tablero(to_integer(11*(yPiezaAct+2) + xPiezaAct)) <= to_unsigned(7,3) when ... else tablero(to_integer(11*(yPiezaAct+2) + xPiezaAct));
  tablero(to_integer(11*(yPiezaAct+1) + (xPiezaAct-1))) <= to_unsigned(7,3) when ... else tablero(to_integer(11*(yPiezaAct+1) + (xPiezaAct-1)));
  
  limpiaTePos2:
  tablero(to_integer(11*yPiezaAct + xPiezaAct)) <= (others => '0') when ... else tablero(to_integer(11*yPiezaAct + xPiezaAct));
  tablero(to_integer(11*yPiezaAct + (xPiezaAct+1))) <= (others => '0') when ... else tablero(to_integer(11*yPiezaAct + (xPiezaAct+1)));
  tablero(to_integer(11*yPiezaAct + (xPiezaAct+2))) <= (others => '0') when ... else tablero(to_integer(11*yPiezaAct + (xPiezaAct+2)));
  tablero(to_integer(11*(yPiezaAct-1) + (xPiezaAct+1))) <= (others => '0') when ... else tablero(to_integer(11*(yPiezaAct-1) + (xPiezaAct+1)));
   
  pintaTePos2:
  tablero(to_integer(11*yPiezaAct + xPiezaAct)) <= to_unsigned(7,3) when ... else tablero(to_integer(11*yPiezaAct + xPiezaAct));
  tablero(to_integer(11*yPiezaAct + (xPiezaAct+1))) <= to_unsigned(7,3) when ... else tablero(to_integer(11*yPiezaAct + (xPiezaAct+1)));
  tablero(to_integer(11*yPiezaAct + (xPiezaAct+2))) <= to_unsigned(7,3) when ... else tablero(to_integer(11*yPiezaAct + (xPiezaAct+2)));
  tablero(to_integer(11*(yPiezaAct-1) + (xPiezaAct+1))) <= to_unsigned(7,3) when ... else tablero(to_integer(11*(yPiezaAct-1) + (xPiezaAct+1)));
  
  limpiaTePos3:
  tablero(to_integer(11*yPiezaAct + xPiezaAct)) <= (others => '0') when ... else tablero(to_integer(11*yPiezaAct + xPiezaAct));
  tablero(to_integer(11*(yPiezaAct+1) + xPiezaAct)) <= (others => '0') when ... else tablero(to_integer(11*(yPiezaAct+1) + xPiezaAct));
  tablero(to_integer(11*(yPiezaAct+2) + xPiezaAct)) <= (others => '0') when ... else tablero(to_integer(11*(yPiezaAct+2) + xPiezaAct));
  tablero(to_integer(11*(yPiezaAct+1) + (xPiezaAct+1))) <= (others => '0') when ... else tablero(to_integer(11*(yPiezaAct+1) + (xPiezaAct+1)));
   
  pintaTePos3:
  tablero(to_integer(11*yPiezaAct + xPiezaAct)) <= to_unsigned(7,3) when ... else tablero(to_integer(11*yPiezaAct + xPiezaAct));
  tablero(to_integer(11*(yPiezaAct+1) + xPiezaAct)) <= to_unsigned(7,3) when ... else tablero(to_integer(11*(yPiezaAct+1) + xPiezaAct));
  tablero(to_integer(11*(yPiezaAct+2) + xPiezaAct)) <= to_unsigned(7,3) when ... else tablero(to_integer(11*(yPiezaAct+2) + xPiezaAct));
  tablero(to_integer(11*(yPiezaAct+1) + (xPiezaAct+1))) <= to_unsigned(7,3) when ... else tablero(to_integer(11*(yPiezaAct+1) + (xPiezaAct+1)));
  
  limpiaTePos4:
  tablero(to_integer(11*yPiezaAct + xPiezaAct)) <= (others => '0') when ... else tablero(to_integer(11*yPiezaAct + xPiezaAct));
  tablero(to_integer(11*yPiezaAct + (xPiezaAct+1))) <= (others => '0') when ... else tablero(to_integer(11*yPiezaAct + (xPiezaAct+1)));
  tablero(to_integer(11*yPiezaAct + (xPiezaAct+2))) <= (others => '0') when ... else tablero(to_integer(11*yPiezaAct + (xPiezaAct+2)));
  tablero(to_integer(11*(yPiezaAct+1) + (xPiezaAct+1))) <= (others => '0') when ... else tablero(to_integer(11*(yPiezaAct+1) + (xPiezaAct+1)));
   
  pintaTePos4:
  tablero(to_integer(11*yPiezaAct + xPiezaAct)) <= to_unsigned(7,3) when ... else tablero(to_integer(11*yPiezaAct + xPiezaAct));
  tablero(to_integer(11*yPiezaAct + (xPiezaAct+1))) <= to_unsigned(7,3) when ... else tablero(to_integer(11*yPiezaAct + (xPiezaAct+1)));
  tablero(to_integer(11*yPiezaAct + (xPiezaAct+2))) <= to_unsigned(7,3) when ... else tablero(to_integer(11*yPiezaAct + (xPiezaAct+2)));
  tablero(to_integer(11*(yPiezaAct+1) + (xPiezaAct+1))) <= to_unsigned(7,3) when ... else tablero(to_integer(11*(yPiezaAct+1) + (xPiezaAct+1)));
  
END syn;
